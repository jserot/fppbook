library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package img_types is
  subtype pixel8 is unsigned(7 downto 0);
end package;

library ieee;
use ieee.std_logic_1164.all;	   
use work.data_types.all;	   

entity tb is
end tb;

architecture struct of tb is

  signal clk: std_logic;
  signal rst: std_logic;
  signal TxWr: std_logic;
  signal TxData: std_logic_vector(7 downto 0);
  signal RxErr: std_logic;
  signal RxRdy: std_logic;
  signal RxData: std_logic_vector(7 downto 0);
  signal TxRdy: std_logic;
  signal RxTx: std_logic;

  constant test_data: int8_array := ( 170, 171, 69 );

begin
  I: entity work.input_tx generic map(test_data) port map(TxWr, TxData, TxRdy);
  T: entity work.tx
    generic map(4, 4)
    port map(clk, TxData, TxWr, TxRdy, RxTx, rst);

  CLOCK: process
  begin
    clk<='1'; wait for 5 ns;
    clk<='0'; wait for 5 ns;
  end process;

  RESET: process
  begin
    rst <= '1'; wait for 5 ns;
    rst <= '0'; wait;
  end process;
end architecture;
